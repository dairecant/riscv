module riscvDemo (

input clk,
input rst,
input [2:0] exControl,
output boot,

);