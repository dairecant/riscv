`timescale 1ns / 1ps
module riscv_imem_tb();

parameter FREQ            = 50000000;
parameter PERIOD          = (1/FREQ)/0.000000001; 
parameter CLK_HALF_PERIOD = PERIOD/2;

parameter INIT_FILE       = "instr_mem_init1.mif";
logic clk_tb,rst_n_tb,en_n_tb,valid_tb;
riscVDat instruction_tb,PC_tb;

riscv_core dut(	
						.clk(clk_tb),
						.rst_n(rst_n_tb),
						.instruction(instruction_tb),
						.pc1(PC_tb),
						.valid(valid_tb)

					);

initial
	begin
		clk_tb = '0;
		forever
			begin
				clk_tb = #(CLK_HALF_PERIOD) ~clk_tb;
			end
	end
					
initial 
	begin
		rst_n_tb = 1'b0;
		#(10*PERIOD) rst_n_tb = 1'b1;
		//$readmemh(INIT_FILE,dut.instr_mem.u0.onchip_memory2_0.the_altsyncram.autogenerated)	;

	
	end
endmodule